* GA CMOS Amp | W=2.628777634427698e-06 L=1e-06 Vbias=1.2225527880022047
.param W=2.628777634427698e-06 L=1e-06 Vbias=1.2225527880022047
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.628777634427698e-06  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 1.2225527880022047 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
