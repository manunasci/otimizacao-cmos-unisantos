* GA CMOS Amp | W=1.0839217174469225e-05 L=1e-06 Vbias=0.8124181163181411
.param W=1.0839217174469225e-05 L=1e-06 Vbias=0.8124181163181411
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.0839217174469225e-05  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.8124181163181411 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
