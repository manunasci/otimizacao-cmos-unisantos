* GA CMOS Amp | W=3.603497878673739e-05 L=9.237339642530373e-07 Vbias=0.5696104521857249
.param W=3.603497878673739e-05 L=9.237339642530373e-07 Vbias=0.5696104521857249
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.603497878673739e-05  L=9.237339642530373e-07
Rload out vdd 10k
Vg  g   0  DC 0.5696104521857249 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
