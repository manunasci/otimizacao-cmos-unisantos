* GA CMOS Amp | W=2.585397349467572e-05 L=2.1461436545397625e-07 Vbias=0.7700576812184586
.param W=2.585397349467572e-05 L=2.1461436545397625e-07 Vbias=0.7700576812184586
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.585397349467572e-05  L=2.1461436545397625e-07
Rload out vdd 10k
Vg  g   0  DC 0.7700576812184586 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
