* GA CMOS Amp | W=1.4006759632267044e-05 L=2.009287462254596e-07 Vbias=1.0147046880768549
.param W=1.4006759632267044e-05 L=2.009287462254596e-07 Vbias=1.0147046880768549
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.4006759632267044e-05  L=2.009287462254596e-07
Rload out vdd 10k
Vg  g   0  DC 1.0147046880768549 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
