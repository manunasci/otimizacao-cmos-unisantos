* GA CMOS Amp | W=1.5726248727690128e-05 L=9.811248163105945e-07 Vbias=0.6213178530783067
.param W=1.5726248727690128e-05 L=9.811248163105945e-07 Vbias=0.6213178530783067
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.5726248727690128e-05  L=9.811248163105945e-07
Rload out vdd 10k
Vg  g   0  DC 0.6213178530783067 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
