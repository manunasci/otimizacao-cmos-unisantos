* GA CMOS Amp | W=4.224271323113583e-05 L=9.084656606712612e-07 Vbias=0.5
.param W=4.224271323113583e-05 L=9.084656606712612e-07 Vbias=0.5
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.224271323113583e-05  L=9.084656606712612e-07
Rload out vdd 10k
Vg  g   0  DC 0.5 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
