* GA CMOS Amp | W=4.2089500969394694e-05 L=3.903627545861094e-07 Vbias=0.5214743958035105
.param W=4.2089500969394694e-05 L=3.903627545861094e-07 Vbias=0.5214743958035105
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.2089500969394694e-05  L=3.903627545861094e-07
Rload out vdd 10k
Vg  g   0  DC 0.5214743958035105 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
