* GA CMOS Amp | W=4.5513078788244845e-05 L=2.3645781825124076e-07 Vbias=0.9578597814576897
.param W=4.5513078788244845e-05 L=2.3645781825124076e-07 Vbias=0.9578597814576897
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.5513078788244845e-05  L=2.3645781825124076e-07
Rload out vdd 10k
Vg  g   0  DC 0.9578597814576897 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
