* GA CMOS Amp | W=7.717802204262605e-06 L=2e-07 Vbias=0.8967406091317973
.param W=7.717802204262605e-06 L=2e-07 Vbias=0.8967406091317973
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=7.717802204262605e-06  L=2e-07
Rload out vdd 10k
Vg  g   0  DC 0.8967406091317973 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
