* GA CMOS Amp | W=2.5505545776505838e-05 L=5.78848012460377e-07 Vbias=0.9045834881909102
.param W=2.5505545776505838e-05 L=5.78848012460377e-07 Vbias=0.9045834881909102
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.5505545776505838e-05  L=5.78848012460377e-07
Rload out vdd 10k
Vg  g   0  DC 0.9045834881909102 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
