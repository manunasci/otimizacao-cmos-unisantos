* GA CMOS Amp | W=3.865758230811834e-05 L=9.98243953993104e-07 Vbias=1.2500833242526772
.param W=3.865758230811834e-05 L=9.98243953993104e-07 Vbias=1.2500833242526772
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.865758230811834e-05  L=9.98243953993104e-07
Rload out vdd 10k
Vg  g   0  DC 1.2500833242526772 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
