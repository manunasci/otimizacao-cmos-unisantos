* GA CMOS Amp | W=2.994731298066147e-05 L=3.66000717742054e-07 Vbias=0.5783697419754558
.param W=2.994731298066147e-05 L=3.66000717742054e-07 Vbias=0.5783697419754558
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.994731298066147e-05  L=3.66000717742054e-07
Rload out vdd 10k
Vg  g   0  DC 0.5783697419754558 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
