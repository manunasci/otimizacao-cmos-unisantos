* GA CMOS Amp | W=2.2207612654295032e-05 L=2.0856037905835396e-07 Vbias=0.742182963358309
.param W=2.2207612654295032e-05 L=2.0856037905835396e-07 Vbias=0.742182963358309
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.2207612654295032e-05  L=2.0856037905835396e-07
Rload out vdd 10k
Vg  g   0  DC 0.742182963358309 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
