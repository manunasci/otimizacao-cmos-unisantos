* GA CMOS Amp | W=4.691708039222585e-05 L=8.266289160596215e-07 Vbias=1.0759767012496233
.param W=4.691708039222585e-05 L=8.266289160596215e-07 Vbias=1.0759767012496233
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.691708039222585e-05  L=8.266289160596215e-07
Rload out vdd 10k
Vg  g   0  DC 1.0759767012496233 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
