* GA CMOS Amp | W=1.9434846082399495e-05 L=1e-06 Vbias=0.578335787156311
.param W=1.9434846082399495e-05 L=1e-06 Vbias=0.578335787156311
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.9434846082399495e-05  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.578335787156311 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
