* GA CMOS Amp | W=8.037292597559787e-06 L=2.0000000000000002e-07 Vbias=1.0698717480125237
.param W=8.037292597559787e-06 L=2.0000000000000002e-07 Vbias=1.0698717480125237
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=8.037292597559787e-06  L=2.0000000000000002e-07
Rload out vdd 10k
Vg  g   0  DC 1.0698717480125237 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
