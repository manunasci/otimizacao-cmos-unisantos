* Amplificador CMOS – W=2.0712752147157204e-05 L=-1.1865744663122963e-08 Vbias=1.0916536908656524
.param W=2.0712752147157204e-05 L=-1.1865744663122963e-08 Vbias=1.0916536908656524

* Biblioteca de processo
.include "C:\Users\holam\OneDrive - Sociedade Visconde de São Leopoldo\Área de Trabalho\otimizacao-cmos-unisantos\cmosedu_models.txt"

* Dispositivo principal (usar modelos 'N' e 'P' do cmosedu_models.txt)
* Aqui usamos apenas um NMOS como exemplo (common-source com carga resistiva)
M1    out in   bias 0   N W=2.0712752147157204e-05 L=-1.1865744663122963e-08
Rload out vdd       10k
Vbias bias 0        DC 1.0916536908656524
Vin   in   0        AC 1
Vdd   vdd  0        DC 1.8

* Análises
.op
.ac dec 100 1 1e9

* Medidas
.measure ac GAIN_LIN  MAX mag(v(out)/v(in))
.measure ac GAIN_DB   MAX db(v(out)/v(in))
* UGBW (unity gain bandwidth) = frequência onde |H(jw)| = 1
.measure ac FC        WHEN mag(v(out)/v(in))=1 CROSS=1
.measure op Idd       FIND I(Vdd)

.end
