* GA CMOS Amp | W=5.204937187065402e-06 L=1e-06 Vbias=0.822111166702319
.param W=5.204937187065402e-06 L=1e-06 Vbias=0.822111166702319
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=5.204937187065402e-06  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.822111166702319 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
