* GA CMOS Amp | W=2.5145720724132312e-05 L=2.0000000000000002e-07 Vbias=1.1973589022736637
.param W=2.5145720724132312e-05 L=2.0000000000000002e-07 Vbias=1.1973589022736637
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.5145720724132312e-05  L=2.0000000000000002e-07
Rload out vdd 10k
Vg  g   0  DC 1.1973589022736637 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
