* GA CMOS Amp | W=8.58703207353758e-06 L=1e-06 Vbias=0.7357224073422363
.param W=8.58703207353758e-06 L=1e-06 Vbias=0.7357224073422363
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=8.58703207353758e-06  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.7357224073422363 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
