* GA CMOS Amp | W=3.080899032084627e-05 L=9.325318427527925e-07 Vbias=0.542510392227586
.param W=3.080899032084627e-05 L=9.325318427527925e-07 Vbias=0.542510392227586
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.080899032084627e-05  L=9.325318427527925e-07
Rload out vdd 10k
Vg  g   0  DC 0.542510392227586 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
