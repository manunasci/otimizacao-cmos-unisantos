* GA CMOS Amp | W=1.53258978432913e-05 L=2.1178509772815867e-07 Vbias=0.6531002292565256
.param W=1.53258978432913e-05 L=2.1178509772815867e-07 Vbias=0.6531002292565256
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.53258978432913e-05  L=2.1178509772815867e-07
Rload out vdd 10k
Vg  g   0  DC 0.6531002292565256 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
