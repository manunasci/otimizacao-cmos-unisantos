* GA CMOS Amp | W=2.886523181248768e-05 L=8.913091852520656e-07 Vbias=0.6004291664758503
.param W=2.886523181248768e-05 L=8.913091852520656e-07 Vbias=0.6004291664758503
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.886523181248768e-05  L=8.913091852520656e-07
Rload out vdd 10k
Vg  g   0  DC 0.6004291664758503 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
