* GA CMOS Amp | W=1.8535638433908004e-06 L=7.427067938629301e-07 Vbias=0.6381294207703707
.param W=1.8535638433908004e-06 L=7.427067938629301e-07 Vbias=0.6381294207703707
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.8535638433908004e-06  L=7.427067938629301e-07
Rload out vdd 10k
Vg  g   0  DC 0.6381294207703707 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
