* Amplificador CMOS � W=7.988850672197389e-06 L=1.834698678492614e-06 Vbias=0.773399127172899
.param W=7.988850672197389e-06 L=1.834698678492614e-06 Vbias=0.773399127172899

* Modelos de fallback
.model nmos NMOS
.model pmos PMOS

* Biblioteca de processo
.include "C:\Users\holam\OneDrive - Sociedade Visconde de S�o Leopoldo\�rea de Trabalho\otimizacao-cmos-unisantos\transistor_model.lib"

* Dispositivos
M1    out in   bias 0   nmos W=7.988850672197389e-06 L=1.834698678492614e-06
Rload out vdd       10k
Vbias bias 0        DC 0.773399127172899
Vin   in   0        AC 1
Vdd   vdd  0        DC 1.8

* An�lises
.op
.ac dec 100 1 1e9

* Medi��es
.measure ac GAIN_LIN MAX mag(v(out)/v(in))
.measure ac GAIN_DB  MAX db(v(out)/v/in))
.measure ac FC       WHEN mag(v(out)/v(in))=GAIN_LIN/sqrt(2)
.measure op  Idd     FIND I(Vdd)

.end
