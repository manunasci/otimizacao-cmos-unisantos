* GA CMOS Amp | W=6.620944666825835e-06 L=6.63809420639884e-07 Vbias=1.0188733071125413
.param W=6.620944666825835e-06 L=6.63809420639884e-07 Vbias=1.0188733071125413
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=6.620944666825835e-06  L=6.63809420639884e-07
Rload out vdd 10k
Vg  g   0  DC 1.0188733071125413 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
