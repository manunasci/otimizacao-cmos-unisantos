* GA CMOS Amp | W=1e-06 L=7.776817081777561e-07 Vbias=0.5
.param W=1e-06 L=7.776817081777561e-07 Vbias=0.5
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1e-06  L=7.776817081777561e-07
Rload out vdd 10k
Vg  g   0  DC 0.5 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
