* GA CMOS Amp | W=1.5787302505900215e-05 L=5.834446853474216e-07 Vbias=1.086873239443484
.param W=1.5787302505900215e-05 L=5.834446853474216e-07 Vbias=1.086873239443484
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.5787302505900215e-05  L=5.834446853474216e-07
Rload out vdd 10k
Vg  g   0  DC 1.086873239443484 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
