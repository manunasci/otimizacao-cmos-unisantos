* GA CMOS Amp | W=4.49390686316207e-06 L=7.115775748802829e-07 Vbias=0.6342616772852195
.param W=4.49390686316207e-06 L=7.115775748802829e-07 Vbias=0.6342616772852195
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.49390686316207e-06  L=7.115775748802829e-07
Rload out vdd 10k
Vg  g   0  DC 0.6342616772852195 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
