* GA CMOS Amp | W=4.54159690306891e-05 L=5.247783701742454e-07 Vbias=0.6230692199139892
.param W=4.54159690306891e-05 L=5.247783701742454e-07 Vbias=0.6230692199139892
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.54159690306891e-05  L=5.247783701742454e-07
Rload out vdd 10k
Vg  g   0  DC 0.6230692199139892 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
