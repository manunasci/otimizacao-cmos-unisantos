* GA CMOS Amp | W=1.3147292602309894e-05 L=2.0000000000000002e-07 Vbias=0.9099795017914397
.param W=1.3147292602309894e-05 L=2.0000000000000002e-07 Vbias=0.9099795017914397
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.3147292602309894e-05  L=2.0000000000000002e-07
Rload out vdd 10k
Vg  g   0  DC 0.9099795017914397 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
