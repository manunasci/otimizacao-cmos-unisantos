* GA CMOS Amp | W=1.3459779271457162e-05 L=2.1190511696978402e-07 Vbias=1.037109541079607
.param W=1.3459779271457162e-05 L=2.1190511696978402e-07 Vbias=1.037109541079607
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.3459779271457162e-05  L=2.1190511696978402e-07
Rload out vdd 10k
Vg  g   0  DC 1.037109541079607 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
