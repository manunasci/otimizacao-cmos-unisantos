* GA CMOS Amp | W=9.859257794762132e-06 L=2.0083754081327224e-07 Vbias=0.5147590137311555
.param W=9.859257794762132e-06 L=2.0083754081327224e-07 Vbias=0.5147590137311555
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=9.859257794762132e-06  L=2.0083754081327224e-07
Rload out vdd 10k
Vg  g   0  DC 0.5147590137311555 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
