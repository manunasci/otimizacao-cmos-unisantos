* GA CMOS Amp | W=1.4644076735765244e-06 L=9.851929830815824e-07 Vbias=0.9778071180199879
.param W=1.4644076735765244e-06 L=9.851929830815824e-07 Vbias=0.9778071180199879
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.4644076735765244e-06  L=9.851929830815824e-07
Rload out vdd 10k
Vg  g   0  DC 0.9778071180199879 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
