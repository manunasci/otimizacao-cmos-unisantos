* GA CMOS Amp | W=4.2754707923220395e-05 L=6.405457320824297e-07 Vbias=0.7584031566436006
.param W=4.2754707923220395e-05 L=6.405457320824297e-07 Vbias=0.7584031566436006
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.2754707923220395e-05  L=6.405457320824297e-07
Rload out vdd 10k
Vg  g   0  DC 0.7584031566436006 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
