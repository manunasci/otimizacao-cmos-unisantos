* GA CMOS Amp | W=9.23408248083964e-06 L=2.1821436450073514e-07 Vbias=1.1605679402867781
.param W=9.23408248083964e-06 L=2.1821436450073514e-07 Vbias=1.1605679402867781
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=9.23408248083964e-06  L=2.1821436450073514e-07
Rload out vdd 10k
Vg  g   0  DC 1.1605679402867781 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
