* GA CMOS Amp | W=7.768493109365587e-06 L=9.852061595991908e-07 Vbias=0.9902726306567183
.param W=7.768493109365587e-06 L=9.852061595991908e-07 Vbias=0.9902726306567183
.options numdgt=6
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=7.768493109365587e-06  L=9.852061595991908e-07
Rload out vdd 10k
Vg  g   0  DC 0.9902726306567183 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 100 1 1e9
.measure ac GAIN_DB  MAX  db(v(out)/v(g))
.measure ac GAIN_LIN MAX  mag(v(out)/v(g))
.measure ac FC WHEN mag(v(out)/v(g))=1 CROSS=1
.measure op Idd param -I(Vdd)
.end
