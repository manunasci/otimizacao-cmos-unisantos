* GA CMOS Amp | W=4.970536543051307e-05 L=5.719529852429772e-07 Vbias=1.1201752930274218
.param W=4.970536543051307e-05 L=5.719529852429772e-07 Vbias=1.1201752930274218
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.970536543051307e-05  L=5.719529852429772e-07
Rload out vdd 10k
Vg  g   0  DC 1.1201752930274218 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
