* GA CMOS Amp | W=1.7875260548570614e-05 L=1e-06 Vbias=0.5890204458474121
.param W=1.7875260548570614e-05 L=1e-06 Vbias=0.5890204458474121
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.7875260548570614e-05  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.5890204458474121 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
