* GA CMOS Amp | W=2.4337293209419226e-05 L=8.417614409410276e-07 Vbias=1.3426985957832667
.param W=2.4337293209419226e-05 L=8.417614409410276e-07 Vbias=1.3426985957832667
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.4337293209419226e-05  L=8.417614409410276e-07
Rload out vdd 10k
Vg  g   0  DC 1.3426985957832667 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
