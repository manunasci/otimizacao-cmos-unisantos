* GA CMOS Amp | W=2.2935766489919234e-05 L=6.888849976093553e-07 Vbias=0.5355635103631733
.param W=2.2935766489919234e-05 L=6.888849976093553e-07 Vbias=0.5355635103631733
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.2935766489919234e-05  L=6.888849976093553e-07
Rload out vdd 10k
Vg  g   0  DC 0.5355635103631733 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
