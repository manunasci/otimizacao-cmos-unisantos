* GA CMOS Amp | W=1e-06 L=8.071499671102273e-07 Vbias=1.1549191672314292
.param W=1e-06 L=8.071499671102273e-07 Vbias=1.1549191672314292
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1e-06  L=8.071499671102273e-07
Rload out vdd 10k
Vg  g   0  DC 1.1549191672314292 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
