* GA CMOS Amp | W=4.191847965103762e-05 L=8.679280041524987e-07 Vbias=1.1965571607027559
.param W=4.191847965103762e-05 L=8.679280041524987e-07 Vbias=1.1965571607027559
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.191847965103762e-05  L=8.679280041524987e-07
Rload out vdd 10k
Vg  g   0  DC 1.1965571607027559 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
