* GA CMOS Amp | W=5.370920977325059e-06 L=7.194236552165659e-07 Vbias=0.5883748446654845
.param W=5.370920977325059e-06 L=7.194236552165659e-07 Vbias=0.5883748446654845
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=5.370920977325059e-06  L=7.194236552165659e-07
Rload out vdd 10k
Vg  g   0  DC 0.5883748446654845 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
