* GA CMOS Amp | W=1.0212118878825219e-05 L=8.572142568151054e-07 Vbias=0.7334855437135861
.param W=1.0212118878825219e-05 L=8.572142568151054e-07 Vbias=0.7334855437135861
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.0212118878825219e-05  L=8.572142568151054e-07
Rload out vdd 10k
Vg  g   0  DC 0.7334855437135861 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
