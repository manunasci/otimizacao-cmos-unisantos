* GA CMOS Amp | W=2.913726687996137e-05 L=5.859410196380134e-07 Vbias=0.543283588422936
.param W=2.913726687996137e-05 L=5.859410196380134e-07 Vbias=0.543283588422936
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.913726687996137e-05  L=5.859410196380134e-07
Rload out vdd 10k
Vg  g   0  DC 0.543283588422936 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
