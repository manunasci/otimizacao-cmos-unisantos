* GA CMOS Amp | W=4.181821040848546e-05 L=8.906362289607569e-07 Vbias=1.0567019733608447
.param W=4.181821040848546e-05 L=8.906362289607569e-07 Vbias=1.0567019733608447
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.181821040848546e-05  L=8.906362289607569e-07
Rload out vdd 10k
Vg  g   0  DC 1.0567019733608447 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
