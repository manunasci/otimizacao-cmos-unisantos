* GA CMOS Amp | W=1.049665674768942e-05 L=3.179704655000608e-07 Vbias=0.8972880288878318
.param W=1.049665674768942e-05 L=3.179704655000608e-07 Vbias=0.8972880288878318
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.049665674768942e-05  L=3.179704655000608e-07
Rload out vdd 10k
Vg  g   0  DC 0.8972880288878318 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
