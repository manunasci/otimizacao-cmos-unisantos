* GA CMOS Amp | W=3.532186634747061e-05 L=6.748079338699678e-07 Vbias=0.7606642335950379
.param W=3.532186634747061e-05 L=6.748079338699678e-07 Vbias=0.7606642335950379
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.532186634747061e-05  L=6.748079338699678e-07
Rload out vdd 10k
Vg  g   0  DC 0.7606642335950379 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
