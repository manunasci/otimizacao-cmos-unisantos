* GA CMOS Amp | W=4.768740289900276e-05 L=4.6783656503563835e-07 Vbias=0.6779066367911027
.param W=4.768740289900276e-05 L=4.6783656503563835e-07 Vbias=0.6779066367911027
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.768740289900276e-05  L=4.6783656503563835e-07
Rload out vdd 10k
Vg  g   0  DC 0.6779066367911027 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
