* GA CMOS Amp | W=3.539196273395511e-05 L=5.259383328528783e-07 Vbias=0.6216269243209289
.param W=3.539196273395511e-05 L=5.259383328528783e-07 Vbias=0.6216269243209289
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.539196273395511e-05  L=5.259383328528783e-07
Rload out vdd 10k
Vg  g   0  DC 0.6216269243209289 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
