* GA CMOS Amp | W=1.5753840922485986e-05 L=6.320155354219852e-07 Vbias=1.0165170473012761
.param W=1.5753840922485986e-05 L=6.320155354219852e-07 Vbias=1.0165170473012761
.options numdgt=6
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.5753840922485986e-05  L=6.320155354219852e-07
Rload out vdd 10k
Vg  g   0  DC 1.0165170473012761 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 100 1 1e9
.measure ac GAIN_DB  MAX  db(v(out)/v(g))
.measure ac GAIN_LIN MAX  mag(v(out)/v(g))
.measure ac FC WHEN mag(v(out)/v(g))=1 CROSS=1
.measure op Idd param -I(Vdd)
.end
