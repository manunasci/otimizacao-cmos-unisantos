* GA CMOS Amp | W=2.8092468391617072e-05 L=6.270842211790859e-07 Vbias=0.6286598305205213
.param W=2.8092468391617072e-05 L=6.270842211790859e-07 Vbias=0.6286598305205213
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.8092468391617072e-05  L=6.270842211790859e-07
Rload out vdd 10k
Vg  g   0  DC 0.6286598305205213 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
