* GA CMOS Amp | W=1.7354183249348018e-05 L=1e-06 Vbias=0.797287200241841
.param W=1.7354183249348018e-05 L=1e-06 Vbias=0.797287200241841
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.7354183249348018e-05  L=1e-06
Rload out vdd 10k
Vg  g   0  DC 0.797287200241841 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
