* GA CMOS Amp | W=1.3829076743266648e-05 L=4.802407805615418e-07 Vbias=0.7229579003982947
.param W=1.3829076743266648e-05 L=4.802407805615418e-07 Vbias=0.7229579003982947
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.3829076743266648e-05  L=4.802407805615418e-07
Rload out vdd 10k
Vg  g   0  DC 0.7229579003982947 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
