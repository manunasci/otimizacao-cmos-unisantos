* GA CMOS Amp | W=4.629461997721569e-05 L=4.444329731807591e-07 Vbias=0.6948286183398787
.param W=4.629461997721569e-05 L=4.444329731807591e-07 Vbias=0.6948286183398787
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.629461997721569e-05  L=4.444329731807591e-07
Rload out vdd 10k
Vg  g   0  DC 0.6948286183398787 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
