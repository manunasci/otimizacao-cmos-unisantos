* GA CMOS Amp | W=9.01890846702332e-06 L=8.964180926543314e-07 Vbias=0.6622431585198771
.param W=9.01890846702332e-06 L=8.964180926543314e-07 Vbias=0.6622431585198771
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=9.01890846702332e-06  L=8.964180926543314e-07
Rload out vdd 10k
Vg  g   0  DC 0.6622431585198771 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
