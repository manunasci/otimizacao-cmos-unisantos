* GA CMOS Amp | W=5.654535879253826e-06 L=2.0729417593674774e-07 Vbias=0.7183596543774623
.param W=5.654535879253826e-06 L=2.0729417593674774e-07 Vbias=0.7183596543774623
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=5.654535879253826e-06  L=2.0729417593674774e-07
Rload out vdd 10k
Vg  g   0  DC 0.7183596543774623 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
