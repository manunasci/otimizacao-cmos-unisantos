* GA CMOS Amp | W=8.143311995923708e-06 L=6.389461675415719e-07 Vbias=0.6439945153000072
.param W=8.143311995923708e-06 L=6.389461675415719e-07 Vbias=0.6439945153000072
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=8.143311995923708e-06  L=6.389461675415719e-07
Rload out vdd 10k
Vg  g   0  DC 0.6439945153000072 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
