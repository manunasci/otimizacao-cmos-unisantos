* GA CMOS Amp | W=9.22759537448246e-06 L=2.0062938479422198e-07 Vbias=1.029784017138696
.param W=9.22759537448246e-06 L=2.0062938479422198e-07 Vbias=1.029784017138696
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=9.22759537448246e-06  L=2.0062938479422198e-07
Rload out vdd 10k
Vg  g   0  DC 1.029784017138696 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
