* GA CMOS Amp | W=2.572244766075149e-05 L=5.715005055775289e-07 Vbias=0.8259307527368991
.param W=2.572244766075149e-05 L=5.715005055775289e-07 Vbias=0.8259307527368991
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.572244766075149e-05  L=5.715005055775289e-07
Rload out vdd 10k
Vg  g   0  DC 0.8259307527368991 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
