* GA CMOS Amp | W=1e-06 L=3.4130810415171946e-07 Vbias=1.432327867956594
.param W=1e-06 L=3.4130810415171946e-07 Vbias=1.432327867956594
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1e-06  L=3.4130810415171946e-07
Rload out vdd 10k
Vg  g   0  DC 1.432327867956594 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
