* GA CMOS Amp | W=3.9446194749976245e-05 L=2.1078099931096333e-07 Vbias=0.8046399740545376
.param W=3.9446194749976245e-05 L=2.1078099931096333e-07 Vbias=0.8046399740545376
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.9446194749976245e-05  L=2.1078099931096333e-07
Rload out vdd 10k
Vg  g   0  DC 0.8046399740545376 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
