* Amplificador CMOS � W=1e-05 L=5e-07 Vbias=0.7
.param W=1e-05 L=5e-07 Vbias=0.7

* Modelos de fallback
.model nmos NMOS
.model pmos PMOS

* Biblioteca de processo
.include "C:\Users\holam\OneDrive - Sociedade Visconde de S�o Leopoldo\�rea de Trabalho\otimizacao-cmos-unisantos\transistor_model.lib"

* Componentes
M1    out in   bias 0   nmos W=1e-05 L=5e-07
Rload out vdd       10k
Vbias bias 0        DC 0.7
Vin   in   0        AC 1
Vdd   vdd  0        DC 1.8

* An�lises
.op
.ac dec 100 1 1e9

* Medi��es no log
.measure ac GMAX MAX mag(v(out)/v(in))
.measure ac FC   WHEN mag(v(out)/v(in))=GMAX/sqrt(2)

.end
