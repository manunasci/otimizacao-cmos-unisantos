* GA CMOS Amp | W=1.0615131066305625e-05 L=2.0422247628166876e-07 Vbias=0.8975232783470165
.param W=1.0615131066305625e-05 L=2.0422247628166876e-07 Vbias=0.8975232783470165
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.0615131066305625e-05  L=2.0422247628166876e-07
Rload out vdd 10k
Vg  g   0  DC 0.8975232783470165 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
