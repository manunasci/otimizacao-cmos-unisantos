* GA CMOS Amp | W=6.251129867681284e-06 L=6.329072896516396e-07 Vbias=0.7376488866317104
.param W=6.251129867681284e-06 L=6.329072896516396e-07 Vbias=0.7376488866317104
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=6.251129867681284e-06  L=6.329072896516396e-07
Rload out vdd 10k
Vg  g   0  DC 0.7376488866317104 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
