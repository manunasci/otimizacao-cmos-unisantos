* GA CMOS Amp | W=8.873223830927035e-06 L=9.723943294255227e-07 Vbias=0.5069468818644127
.param W=8.873223830927035e-06 L=9.723943294255227e-07 Vbias=0.5069468818644127
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=8.873223830927035e-06  L=9.723943294255227e-07
Rload out vdd 10k
Vg  g   0  DC 0.5069468818644127 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
