* GA CMOS Amp | W=3.5174662158511296e-05 L=5.23424933237009e-07 Vbias=1.4721947321711004
.param W=3.5174662158511296e-05 L=5.23424933237009e-07 Vbias=1.4721947321711004
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.5174662158511296e-05  L=5.23424933237009e-07
Rload out vdd 10k
Vg  g   0  DC 1.4721947321711004 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
