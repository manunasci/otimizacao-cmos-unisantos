* GA CMOS Amp | W=4.430009205494142e-05 L=9.526119679626481e-07 Vbias=1.3056357081452707
.param W=4.430009205494142e-05 L=9.526119679626481e-07 Vbias=1.3056357081452707
.options numdgt=6
.include "models.lib"
* Device
M1  out g  0  0  N  W=4.430009205494142e-05  L=9.526119679626481e-07
Rload out vdd 10k
Vg  g   0  DC 1.3056357081452707 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 100 1 1e9
.measure ac GAIN_DB  MAX  db(v(out)/v(g))
.measure ac GAIN_LIN MAX  mag(v(out)/v(g))
.measure ac FC WHEN mag(v(out)/v(g))=1 CROSS=1
.measure op Idd FIND I(Vdd)
.end
