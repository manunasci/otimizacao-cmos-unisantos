* GA CMOS Amp | W=1.5379070469543866e-05 L=9.783637611803528e-07 Vbias=0.8406286737807008
.param W=1.5379070469543866e-05 L=9.783637611803528e-07 Vbias=0.8406286737807008
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.5379070469543866e-05  L=9.783637611803528e-07
Rload out vdd 10k
Vg  g   0  DC 0.8406286737807008 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
