* GA CMOS Amp | W=2.2931630592261437e-05 L=4.985692553771025e-07 Vbias=0.5873381740588752
.param W=2.2931630592261437e-05 L=4.985692553771025e-07 Vbias=0.5873381740588752
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=2.2931630592261437e-05  L=4.985692553771025e-07
Rload out vdd 10k
Vg  g   0  DC 0.5873381740588752 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
