* Amplificador CMOS - W=4.070484377450471e-05 L=7.601026610045998e-07 Vbias=1.466084216534019
.param W=4.070484377450471e-05 L=7.601026610045998e-07 Vbias=1.466084216534019

* Modelos de fallback
.model nmos NMOS
.model pmos PMOS

* Biblioteca de processo
.include "C:\Users\holam\OneDrive - Sociedade Visconde de S�o Leopoldo\�rea de Trabalho\otimizacao-cmos-unisantos\transistor_model.lib"

* Dispositivos
M1    out in   bias 0   nmos W=4.070484377450471e-05 L=7.601026610045998e-07
Rload out vdd       10k
Vbias bias 0        DC 1.466084216534019
Vin   in   0        AC 1
Vdd   vdd  0        DC 1.8

* An�lises
.op
.ac dec 100 1 1e9

* Medi��es
.measure ac GAIN_LIN MAX mag(v(out)/v(in))
.measure ac GAIN_DB  MAX db(v(out)/v(in))
.measure ac FC       WHEN mag(v(out)/v(in))=GAIN_LIN/sqrt(2)
.measure op  Idd     FIND I(Vdd)

.end
