* GA CMOS Amp | W=5e-05 L=2.096397733682079e-07 Vbias=0.810035335418613
.param W=5e-05 L=2.096397733682079e-07 Vbias=0.810035335418613
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=5e-05  L=2.096397733682079e-07
Rload out vdd 10k
Vg  g   0  DC 0.810035335418613 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
