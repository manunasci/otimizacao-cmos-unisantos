* GA CMOS Amp | W=3.974698015793619e-05 L=3.4018036538324214e-07 Vbias=1.4457714277153724
.param W=3.974698015793619e-05 L=3.4018036538324214e-07 Vbias=1.4457714277153724
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=3.974698015793619e-05  L=3.4018036538324214e-07
Rload out vdd 10k
Vg  g   0  DC 1.4457714277153724 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
