* GA CMOS Amp | W=1.7961368287577085e-06 L=9.900908579105005e-07 Vbias=1.218738405366215
.param W=1.7961368287577085e-06 L=9.900908579105005e-07 Vbias=1.218738405366215
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=1.7961368287577085e-06  L=9.900908579105005e-07
Rload out vdd 10k
Vg  g   0  DC 1.218738405366215 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 400 1 1e9
.save V(out)
.end
