* GA CMOS Amp | W=4.352921277097167e-05 L=9.902986468048787e-07 Vbias=1.1384501006760075
.param W=4.352921277097167e-05 L=9.902986468048787e-07 Vbias=1.1384501006760075
.options numdgt=6
.options plotwinsize=0
.include "models.lib"
* Device
M1  out g  0  0  N_1u  W=4.352921277097167e-05  L=9.902986468048787e-07
Rload out vdd 10k
Vg  g   0  DC 1.1384501006760075 AC 1
Vdd vdd 0  DC 1.8
.op
.ac dec 200 1 1e9
.save V(out) V(g)
.end
